entity stopwatch is
end entity stopwatch;

architecture structural of stopwatch is

begin

end architecture structural;
